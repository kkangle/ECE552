module ALU_tb()