module BitCell(clk, rst, D, WriteEnable, ReadEnable1, ReadEnable2, Bitline1, Bitline2);

input clk,  
input rst, 
input D, 
input WriteEnable, 
input ReadEnable1, 
input ReadEnable2, 
inout Bitline1, 
inout Bitline2



endmodule
